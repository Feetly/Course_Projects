bjt bias 3

.include /home/student/student/Documents/bjt/QN2222.txt
vbb 1 0 dc 15v
r1 1 2 100
q1 3 2 4 Q2N2222A 
r2 2 0 100
r3 5 3 100
r4 4 0 100
v5 6 0 dc 5
vd 6 5 dc 0

.control
dc vbb 0 20 0.2 
run

plot vd#branch vs v(2)
print vd#branch v(2)
.endc
.END
