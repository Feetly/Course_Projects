I-V Characteristics of CD4007
*Including the CD4007 model file
.include /home/student/student/Documents/nmos/cd4007.txt
vgs 1 0 dc 5v
*Specifying NMOS in this manner-
*name drain gate source body modelname as in model file
m1 2 1 0 0 MN4007 
*DC source of 0v to measure current
vid 3 2 dc 0v
vdd 3 0 dc 5v

.control
dc vdd 0 5 .1 vgs 0 5 1 
run
plot vid#branch  xlabel 'Vds' ylabel 'Ids' title 'V-I Characteristics'
print vid#branch v(2)
.endc
.end
